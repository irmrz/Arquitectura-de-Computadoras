module execute (input logic 			 AluSrc,
					 input logic [3:0]    AluControl,
					 input logic [63:0]	 PC_E,
												 signlmm_E,
												 readData1_E,
												 readData2_E,
					 output logic [63:0]  PCBranch_E,
												 aluResult_E,
												 writeData_E,
					 output logic 			 zero_E);

	
endmodule					 